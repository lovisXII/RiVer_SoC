library ieee; 
use ieee.std_logic_1164.all;

package util is 
    constant kernel_adr : std_logic_vector(31 downto 0) := x"F0000000"; 
    constant one_ext_32 : std_logic_vector(31 downto 0) := x"00000001"; 
end util; 

package body util is 
    
end util; 