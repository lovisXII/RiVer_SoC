library ieee; 
use ieee.std_logic_1164.all;

package util is 
    constant kernel_adr : std_logic_vector(31 downto 0) := x"80000000"; 

end util; 

package body util is 
    
end util; 